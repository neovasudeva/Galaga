// user_ship.sv
// used to control the movement of user_ship
// also gives control signals to color_mapper.sv for drawing



module  user_ship ( input         Clk,           // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
					input [7:0]	  keycode,				 // pass key pressed into user_ship.sv
					output 		  is_user_ship,		 // whether current drawing pixel is the user_ship
					output [23:0] user_ship_data,		 // sends color of user ship
					output [9:0]  x_pos,
					output [9:0]  y_pos
              );
    
    parameter [9:0] User_Ship_X_Center = 10'd320;  // Center position on the X axis
    parameter [9:0] User_Ship_Y_Center = 10'd240;  // Center position on the Y axis
    parameter [9:0] User_Ship_X_Min = 10'd0;       // Leftmost point on the X axis
    parameter [9:0] User_Ship_X_Max = 10'd639;     // Rightmost point on the X axis
    parameter [9:0] User_Ship_Y_Min = 10'd0;       // Topmost point on the Y axis
    parameter [9:0] User_Ship_Y_Max = 10'd479;     // Bottommost point on the Y axis
    parameter [9:0] User_Ship_X_Step = 10'd1;      // Step size on the X axis
    parameter [9:0] User_Ship_Y_Step = 10'd1;      // Step size on the Y axis
    parameter [9:0] User_Ship_Size = 10'd40;       // User_Ship's size (40x40)
    
    logic [9:0] User_Ship_X_Motion, User_Ship_Y_Motion, User_Ship_X_Pos, User_Ship_Y_Pos;
    logic [9:0] User_Ship_X_Pos_in, User_Ship_X_Motion_in, User_Ship_Y_Pos_in, User_Ship_Y_Motion_in;
	 
	 assign x_pos = User_Ship_X_Pos;
	 assign y_pos = User_Ship_Y_Pos;
    
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    // Update registers
    always_ff @ (posedge Clk)
    begin
        if (Reset)
        begin
            User_Ship_X_Pos <= User_Ship_X_Center;
            User_Ship_Y_Pos <= User_Ship_Y_Max - User_Ship_Size;	// start at the bottom
            User_Ship_X_Motion <= User_Ship_X_Step;
            User_Ship_Y_Motion <= 10'd0; //User_Ship_Y_Step;
        end
        else
        begin
            User_Ship_X_Pos <= User_Ship_X_Pos_in;
            User_Ship_Y_Pos <= User_Ship_Y_Pos_in;
            User_Ship_X_Motion <= User_Ship_X_Motion_in;
            User_Ship_Y_Motion <= User_Ship_Y_Motion_in;
        end
    end
    //////// Do not modify the always_ff blocks. ////////
    
    // You need to modify always_comb block.
    always_comb
    begin
        // By default, keep motion and position unchanged
        User_Ship_X_Pos_in = User_Ship_X_Pos;
        User_Ship_Y_Pos_in = User_Ship_Y_Pos;
        User_Ship_X_Motion_in = User_Ship_X_Motion;
        User_Ship_Y_Motion_in = User_Ship_Y_Motion;
        
        // Update position and motion only at rising edge of frame clock
        if (frame_clk_rising_edge)
        begin
            // Be careful when using comparators with "logic" datatype because compiler treats 
            //   both sides of the operator as UNSIGNED numbers.
            // e.g. User_Ship_Y_Pos - Ball_Size <= User_Ship_Y_Min 
            // If User_Ship_Y_Pos is 0, then User_Ship_Y_Pos - Ball_Size will not be -4, but rather a large positive number.
				
				// handle keys -> only go left and right
				unique case(keycode)
					8'h04: begin			// A -> go left
						User_Ship_Y_Motion_in = 10'd0;
						User_Ship_X_Motion_in = (~(User_Ship_X_Step) + 1'b1);
					end
					8'h07: begin			// D -> go right
						User_Ship_Y_Motion_in = 10'd0;
						User_Ship_X_Motion_in = User_Ship_X_Step;
					end
					default: begin			// maintain current heading if no keys are pressed
						User_Ship_X_Motion_in = User_Ship_X_Motion;
						User_Ship_Y_Motion_in = User_Ship_Y_Motion;
					end
				endcase
					
				// handle edges -> left and right edges
				if (User_Ship_X_Pos + User_Ship_Size >= User_Ship_X_Max) begin // Ball is at right edge, BOUNCE!
					 User_Ship_X_Motion_in = (~(User_Ship_Y_Step) + 1'b1);
					 User_Ship_Y_Motion_in = 10'd0;
				end
				else if (User_Ship_X_Pos <= User_Ship_X_Min + User_Ship_Size)	begin // Ball is at left edge, BOUNCE!
					 User_Ship_X_Motion_in = User_Ship_X_Step;
					 User_Ship_Y_Motion_in = 10'd0;
				end
        
            // Update the ball's position with its motion
            User_Ship_X_Pos_in = User_Ship_X_Pos + User_Ship_X_Motion;
            User_Ship_Y_Pos_in = User_Ship_Y_Pos + User_Ship_Y_Motion;
        end
    end
	 
	     // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
	 
	 logic [10:0] user_ship_addr;
    always_comb begin
        if ( DrawX >= User_Ship_X_Pos && DrawX < User_Ship_X_Pos + User_Ship_Size &&
				DrawY >= User_Ship_Y_Pos && DrawY < User_Ship_Y_Pos + User_Ship_Size ) begin
				user_ship_addr = (DrawY - User_Ship_Y_Pos) * User_Ship_Size + (DrawX - User_Ship_X_Pos);
				// don't color in background of ship
				if (user_ship_data == 24'h002000) 
					is_user_ship = 1'b0;
				else
					is_user_ship = 1'b1;
		  end
        else begin
				user_ship_addr = 11'h00;	// match background
            is_user_ship = 1'b0;
		  end
    end
	 
	 // get color data of user_ship via on chip memory
	 shipRAM sr(.read_address (user_ship_addr), .Clk (Clk), .data_out(user_ship_data) );
    
endmodule