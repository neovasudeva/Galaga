// sprite roms
// i hope i have enough memory for this garbo


// galaga logo
module galaga_rom (input [3:0] addr,
						output [95:0] data);

	// rom stuff
	logic [0:15][95:0] ROM;
	assign ROM = {
		
		// Galaga
		96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000011111111000000000011000000001111111100000000000000110000000000001111111100000000001100000000,  
      96'b001111000011110000001111110000000011110000000000000011111100000000111100001111000000111111000000,  
      96'b111100000000110000111100111100000011110000000000001111001111000011110000000011000011110011110000,  
      96'b111100000000000011110000001111000011110000000000111100000011110011110000000000001111000000111100,  
      96'b111100000000000011110000001111000011110000000000111100000011110011110000000000001111000000111100,  
      96'b111100111111110011111111111111000011110000000000111111111111110011110011111111001111111111111100,  
      96'b111100000011110011110000001111000011110000000000111100000011110011110000001111001111000000111100,  
      96'b111100000011110011110000001111000011110000000000111100000011110011110000001111001111000000111100,  
      96'b001111000011110011110000001111000011110000001100111100000011110000111100001111001111000000111100,  
      96'b000011111100110011110000001111001111111111111100111100000011110000001111110011001111000000111100,  
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
		
	};
	
	assign data[95:0] = ROM[addr];
		
endmodule		



// game over logo
module gameover_rom (input [3:0] addr,
						output [127:0] data);

	// rom stuff
	logic [0:15][127:0] ROM;
	assign ROM = {
		
		// Gameover
		128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      128'b00001111111100000000001100000000111100000000111111111111111111000011111111110000111100000000111111111111111111001111111111110000,  
      128'b00111100001111000000111111000000111111000011111100111100001111001111000000111100111100000000111100111100001111000011110000111100,  
      128'b11110000000011000011110011110000111111111111111100111100000011001111000000111100111100000000111100111100000011000011110000111100,  
      128'b11110000000000001111000000111100111111111111111100111100110000001111000000111100111100000000111100111100110000000011110000111100,  
      128'b11110000000000001111000000111100111100111100111100111111110000001111000000111100111100000000111100111111110000000011111111110000,  
      128'b11110011111111001111111111111100111100000000111100111100110000001111000000111100111100000000111100111100110000000011110000111100,  
      128'b11110000001111001111000000111100111100000000111100111100000000001111000000111100111100000000111100111100000000000011110000111100,  
      128'b11110000001111001111000000111100111100000000111100111100000011001111000000111100001111000011110000111100000011000011110000111100,  
      128'b00111100001111001111000000111100111100000000111100111111001111001111000000111100000011111111000000111111001111000011110000111100,  
      128'b00001111110011001111000000111100111100000000111111111111111111000011111111110000000000111100000011111111111111001111110000111110,  
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

	};
	
	assign data[127:0] = ROM[addr];
		
endmodule		


// press enter logo
module press_start_rom (input [2:0] addr,
								output [54:0] data);
								
	// rom stuff
	logic [0:4][54:0] ROM;
	assign ROM = {
		
		// Press enter
		55'b1111011100111100111001110000001111010001111111111011100,
		55'b1001010010100001000010000000001000011001001001000010010,
		55'b1111011100111000111001110000001110010101001001110011100,
		55'b1000010100100000000100001000001000010011001001000010100,
		55'b1000010010111100111001110000001111010001001001111010010
		
	};
	
	assign data[54:0] = ROM[addr];
	
endmodule





// you win logo
module you_win_rom (input [3:0] addr,
						output [111:0] data);

	// rom stuff
	logic [0:15][111:0] ROM;
	assign ROM = {
		
		// Galaga
		112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      112'b1111000000001110100111111111100011110000000011110000000000000000111100000000111100001111111100001111000000111100,  
      112'b1111000000001110111110000001111011110000000011110000000000000000111100000000111100000011110000001111110000111100,  
      112'b1111000000001110111110000001111011110000000011110000000000000000111100000000111100000011110000001111111000111100,  
      112'b0011110000111100011110000001111011110000000011110000000000000000111100000000111100000011110000001111111111111100,  
      112'b0000111111110000011110000001111011110000000011110000000000000000111100011000111100000011110000001111001111111100,  
      112'b0000001111000000011110000001111011110000000011110000000000000000111100111100111100000011110000001111000011111100,  
      112'b0000001111000000011110000001111011110000000011110000000000000000111111111111111100000011110000001111000000111100,  
      112'b0000001111000000011110000001111001111000000111100000000000000000111111111111111100000011110000001111000000111100,  
      112'b0000001111000000011110000001111000111111111111000000000000000000111111000011111100000011110000001111000000111100,  
      112'b0000111111110000000111111111100000001111111100000000000000000000111100000000111100001111111100001111000000111100,  
      112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
		
	};
	
	assign data[111:0] = ROM[addr];
		
endmodule		
