// sprite roms
// i hope i have enough memory for this garbo


// galaga logo
module galaga_rom (input [3:0] addr,
						output [95:0] data);

	// rom stuff
	logic [0:15][95:0] ROM;
	assign ROM = {
		
		// G
		96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000011111111000000000011000000001111111100000000000000110000000000001111111100000000001100000000,  
      96'b001111000011110000001111110000000011110000000000000011111100000000111100001111000000111111000000,  
      96'b111100000000110000111100111100000011110000000000001111001111000011110000000011000011110011110000,  
      96'b111100000000000011110000001111000011110000000000111100000011110011110000000000001111000000111100,  
      96'b111100000000000011110000001111000011110000000000111100000011110011110000000000001111000000111100,  
      96'b111100111111110011111111111111000011110000000000111111111111110011110011111111001111111111111100,  
      96'b111100000011110011110000001111000011110000000000111100000011110011110000001111001111000000111100,  
      96'b111100000011110011110000001111000011110000000000111100000011110011110000001111001111000000111100,  
      96'b001111000011110011110000001111000011110000001100111100000011110000111100001111001111000000111100,  
      96'b000011111100110011110000001111001111111111111100111100000011110000001111110011001111000000111100,  
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
		
	};
	
	assign data[95:0] = ROM[addr];
		
endmodule		



// game over logo
module gameover_rom (input [3:0] addr,
						output [127:0] data);

	// rom stuff
	logic [0:15][0:127] ROM;
	assign ROM = {
		
		// G
		96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b00001111111100000000001100000000111100000000111111111111111111000011111111110000111100000000111111111111111111001111111111110000,  
      96'b00111100001111000000111111000000111111000011111100111100001111001111000000111100111100000000111100111100001111000011110000111100,  
      96'b11110000000011000011110011110000111111111111111100111100000011001111000000111100111100000000111100111100000011000011110000111100,  
      96'b11110000000000001111000000111100111111111111111100111100110000001111000000111100111100000000111100111100110000000011110000111100,  
      96'b11110000000000001111000000111100111100111100111100111111110000001111000000111100111100000000111100111111110000000011111111110000,  
      96'b11110011111111001111111111111100111100000000111100111100110000001111000000111100111100000000111100111100110000000011110000111100,  
      96'b11110000001111001111000000111100111100000000111100111100000000001111000000111100111100000000111100111100000000000011110000111100,  
      96'b11110000001111001111000000111100111100000000111100111100000011001111000000111100001111000011110000111100000011000011110000111100,  
      96'b00111100001111001111000000111100111100000000111100111111001111001111000000111100000011111111000000111111001111000011110000111100,  
      96'b00001111110011001111000000111100111100000000111111111111111111000011111111110000000000111100000011111111111111001111110000111110,  
      96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 
      96'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

	};
	
	assign data = ROM[addr];
		
endmodule		
